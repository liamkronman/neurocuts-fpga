
package tree_constants;
    parameter TOTAL_NODES = 50251;
    parameter TOTAL_RULES = 40348;
    parameter MAX_CHILDREN_PER_NODE = 32;
    parameter MAX_RULES_PER_NODE = 16;
endpackage
