
package tree_constants;
    parameter TOTAL_NODES = 24997;
    parameter TOTAL_RULES = 22788;
    parameter MAX_CHILDREN_PER_NODE = 32;
    parameter MAX_RULES_PER_NODE = 16;
endpackage
