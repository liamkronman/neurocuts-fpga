
module neuro_cuts(
    input logic[1:0] a,
    output logic b
);
    assign b = a;
endmodule : neuro_cuts