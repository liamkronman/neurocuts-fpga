

module node(
    logic does_partition,
    rule_s rule
);

endmodule