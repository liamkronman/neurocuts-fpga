
package tree_constants;
    parameter TOTAL_NODES = 370;
    parameter TOTAL_RULES = 317;
    parameter MAX_CHILDREN_PER_NODE = 17;
    parameter MAX_RULES_PER_NODE = 16;
endpackage
